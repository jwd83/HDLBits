/*

Implement the following circuit:

*/

module top_module (
    input clk,
    input resetn,   // synchronous reset
    input in,
    output out);

endmodule
