// A "population count" circuit counts the number of '1's in an input vector.
// Build a population count circuit for a 255-bit input vector.


module top_module(
    input [254:0] in,
    output [7:0] out );

endmodule
